module SNN_Core(

);
endmodule