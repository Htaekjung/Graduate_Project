module CNN_Core(

);
endmodule